// Casey Silcox
// August Avantaggio
// EE 371
// Lab 5
// This program
module DE1_SoC(CLOCK_50, KEY, SW, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0, GPIO_0);

	
endmodule
